module top (input i, output o, input clk);
	assign o = i;
endmodule
