module top (input i, output o, input rce);
	assign o = i;
endmodule
